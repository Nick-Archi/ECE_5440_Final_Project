/* 	Module: CheckMemory
*
* 	Description: Takes the user’s ID and checks the memory in order to access the user’s specified level 
* (if not a guest) and high score. (RAM/ROM)
*
*	Created By: Nicholas
*
*/

module CheckMemory(password, displayLevel);






endmodule
