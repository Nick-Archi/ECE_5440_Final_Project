/* 	Module: UserLogin
* 	Description: Takes the user’s inputted password and 
*	sends this 4 digit value to the CheckMemory module.
*
*	Created By: Nicholas
*
*/

module UserLogin();



endmodule